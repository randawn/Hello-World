
class axi_seq_item extends uvm_sequence_item;
    `uvm_object_utils(axi_seq_item)


endclass: axi_seq_item

