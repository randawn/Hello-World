module t0;
t1 t1(.*);
t2 t2(.*);
endmodule
