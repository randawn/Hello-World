module t2(
    input a,
    output b
);
endmodule
