module t1(
    output a,
    input b
);
endmodule
